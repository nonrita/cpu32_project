`timescale 1ns/1ps

module xor32 (
    input  wire [31:0] A,
    input  wire [31:0] B,
    output wire [31:0] Y
);
    assign Y = A ^ B;
endmodule
